
`timescale 1ns/1ps
module Stage1 (
    input  a,
    input  b,
    output  c
);

    assign c= a & b;

    
endmodule