`timescale 1ns/1ps
module ForReplica #(
    parameter N =4 ;
) (
    
);
    
endmodule